library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity charmem is
  port (clk:  in std_logic;
		  row1: in  std_logic_vector(5 downto 0); -- row address for display side
		  col1: in  std_logic_vector(6 downto 0); -- column address for display
		  out1: out std_logic_vector(6 downto 0); -- character to be displayed
		  row2: in  std_logic_vector(5 downto 0); -- row address for input
		  col2: in  std_logic_vector(6 downto 0); -- column address for input
		  in2:  in  std_logic_vector(6 downto 0); -- character to be input
		  writec: in std_logic; -- write one char (int2) at row2,col2
		  clear:  in std_logic; -- clear the screen (memory)
		  scroll: in std_logic); -- scroll the screen (memory)
end charmem;

architecture behavioral of charmem is
  type char_ram_type is array (0 to 8191) of integer range 0 to 127;
  signal char_ram: char_ram_type := (
62,32,73,102,32,119,101,32,97,114,101,32,109,97,114,107,39,100,32,116,111,32,100,
105,101,44,32,119,101,32,97,114,101,32,101,110,111,119,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,
32,84,111,32,100,111,32,111,117,114,32,99,111,117,110,116,114,121,32,108,111,115,
115,59,32,97,110,100,32,105,102,32,116,111,32,108,105,118,101,44,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,62,32,84,104,101,32,102,101,119,101,114,32,109,101,110,44,32,116,104,101,32,103,
114,101,97,116,101,114,32,115,104,97,114,101,32,111,102,32,104,111,110,111,117,
114,46,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,62,32,71,111,100,39,115,32,119,105,108,108,33,32,73,32,112,114,
97,121,32,116,104,101,101,44,32,119,105,115,104,32,110,111,116,32,111,110,101,32,
109,97,110,32,109,111,114,101,46,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,66,121,32,74,111,118,101,44,32,73,32,97,
109,32,110,111,116,32,99,111,118,101,116,111,117,115,32,102,111,114,32,103,111,
108,100,44,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,78,111,114,32,99,97,114,101,32,73,32,119,
104,111,32,100,111,116,104,32,102,101,101,100,32,117,112,111,110,32,109,121,32,
99,111,115,116,59,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,73,116,32,121,101,97,114,110,115,32,109,
101,32,110,111,116,32,105,102,32,109,101,110,32,109,121,32,103,97,114,109,101,110,
116,115,32,119,101,97,114,59,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,83,117,99,104,32,111,117,116,119,
97,114,100,32,116,104,105,110,103,115,32,100,119,101,108,108,32,110,111,116,32,
105,110,32,109,121,32,100,101,115,105,114,101,115,46,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,66,117,116,32,
105,102,32,105,116,32,98,101,32,97,32,115,105,110,32,116,111,32,99,111,118,101,
116,32,104,111,110,111,117,114,44,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,73,32,97,109,32,
116,104,101,32,109,111,115,116,32,111,102,102,101,110,100,105,110,103,32,115,111,
117,108,32,97,108,105,118,101,46,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,78,111,44,32,102,
97,105,116,104,44,32,109,121,32,99,111,122,44,32,119,105,115,104,32,110,111,116,
32,97,32,109,97,110,32,102,114,111,109,32,69,110,103,108,97,110,100,46,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,71,
111,100,39,115,32,112,101,97,99,101,33,32,73,32,119,111,117,108,100,32,110,111,
116,32,108,111,115,101,32,115,111,32,103,114,101,97,116,32,97,110,32,104,111,110,
111,117,114,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,62,32,65,115,32,111,110,101,32,109,97,110,32,109,111,114,101,32,109,101,
116,104,105,110,107,115,32,119,111,117,108,100,32,115,104,97,114,101,32,102,114,
111,109,32,109,101,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,70,111,114,32,116,104,101,32,98,101,115,116,32,
104,111,112,101,32,73,32,104,97,118,101,46,32,79,44,32,100,111,32,110,111,116,32,
119,105,115,104,32,111,110,101,32,109,111,114,101,33,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,82,97,116,104,101,114,32,
112,114,111,99,108,97,105,109,32,105,116,44,32,87,101,115,116,109,111,114,101,108,
97,110,100,44,32,116,104,114,111,117,103,104,32,109,121,32,104,111,115,116,44,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,84,
104,97,116,32,104,101,32,119,104,105,99,104,32,104,97,116,104,32,110,111,32,115,
116,111,109,97,99,104,32,116,111,32,116,104,105,115,32,102,105,103,104,116,44,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,62,32,76,101,116,32,104,105,109,32,100,101,112,97,114,116,59,32,104,105,115,
32,112,97,115,115,112,111,114,116,32,115,104,97,108,108,32,98,101,32,109,97,100,
101,44,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,62,32,65,110,100,32,99,114,111,119,110,115,32,102,111,114,32,99,
111,110,118,111,121,32,112,117,116,32,105,110,116,111,32,104,105,115,32,112,117,
114,115,101,59,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,87,101,32,119,111,117,108,100,32,110,111,116,
32,100,105,101,32,105,110,32,116,104,97,116,32,109,97,110,39,115,32,99,111,109,
112,97,110,121,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,84,104,97,116,32,102,101,97,114,115,32,
104,105,115,32,102,101,108,108,111,119,115,104,105,112,32,116,111,32,100,105,101,
32,119,105,116,104,32,117,115,46,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,84,104,105,115,32,100,97,121,
32,105,115,32,99,97,108,108,39,100,32,116,104,101,32,102,101,97,115,116,32,111,
102,32,67,114,105,115,112,105,97,110,46,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,72,101,32,116,104,97,
116,32,111,117,116,108,105,118,101,115,32,116,104,105,115,32,100,97,121,44,32,97,
110,100,32,99,111,109,101,115,32,115,97,102,101,32,104,111,109,101,44,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,87,
105,108,108,32,115,116,97,110,100,32,97,32,116,105,112,45,116,111,101,32,119,104,
101,110,32,116,104,105,115,32,100,97,121,32,105,115,32,110,97,109,39,100,44,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,62,32,65,110,100,32,114,111,117,115,101,32,104,105,109,32,97,116,32,116,104,101,
32,110,97,109,101,32,111,102,32,67,114,105,115,112,105,97,110,46,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,62,32,72,101,32,116,104,97,116,32,115,104,97,108,108,32,108,105,118,101,32,
116,104,105,115,32,100,97,121,44,32,97,110,100,32,115,101,101,32,111,108,100,32,
97,103,101,44,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,62,32,87,105,108,108,32,121,101,97,114,108,121,32,111,110,32,
116,104,101,32,118,105,103,105,108,32,102,101,97,115,116,32,104,105,115,32,110,
101,105,103,104,98,111,117,114,115,44,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,65,110,100,32,115,97,121,32,34,84,
111,45,109,111,114,114,111,119,32,105,115,32,83,97,105,110,116,32,67,114,105,115,
112,105,97,110,46,34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,84,104,101,110,32,119,105,108,108,
32,104,101,32,115,116,114,105,112,32,104,105,115,32,115,108,101,101,118,101,32,
97,110,100,32,115,104,111,119,32,104,105,115,32,115,99,97,114,115,44,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,65,110,
100,32,115,97,121,32,34,84,104,101,115,101,32,119,111,117,110,100,115,32,73,32,
104,97,100,32,111,110,32,67,114,105,115,112,105,97,110,39,115,32,100,97,121,46,
34,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,62,32,79,108,100,32,109,101,110,32,102,111,114,103,101,116,59,32,121,101,116,
32,97,108,108,32,115,104,97,108,108,32,98,101,32,102,111,114,103,111,116,44,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,62,32,66,117,116,32,104,101,39,108,108,32,114,101,109,101,109,98,101,
114,44,32,119,105,116,104,32,97,100,118,97,110,116,97,103,101,115,44,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,62,32,87,104,97,116,32,102,101,97,116,115,32,104,101,32,100,105,100,
32,116,104,97,116,32,100,97,121,46,32,84,104,101,110,32,115,104,97,108,108,32,111,
117,114,32,110,97,109,101,115,44,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,70,97,109,105,108,105,97,114,32,105,110,32,
104,105,115,32,109,111,117,116,104,32,97,115,32,104,111,117,115,101,104,111,108,
100,32,119,111,114,100,115,45,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,72,97,114,114,121,32,116,104,101,
32,75,105,110,103,44,32,66,101,100,102,111,114,100,32,97,110,100,32,69,120,101,
116,101,114,44,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,87,97,114,119,105,99,107,32,97,110,
100,32,84,97,108,98,111,116,44,32,83,97,108,105,115,98,117,114,121,32,97,110,100,
32,71,108,111,117,99,101,115,116,101,114,45,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,66,101,32,105,110,32,116,
104,101,105,114,32,102,108,111,119,105,110,103,32,99,117,112,115,32,102,114,101,
115,104,108,121,32,114,101,109,101,109,98,39,114,101,100,46,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,84,104,
105,115,32,115,116,111,114,121,32,115,104,97,108,108,32,116,104,101,32,103,111,
111,100,32,109,97,110,32,116,101,97,99,104,32,104,105,115,32,115,111,110,59,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,62,32,65,110,100,32,67,114,105,115,112,105,110,32,67,114,105,115,112,105,97,110,
32,115,104,97,108,108,32,110,101,39,101,114,32,103,111,32,98,121,44,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,62,32,70,114,111,109,32,116,104,105,115,32,100,97,121,32,116,111,32,116,104,
101,32,101,110,100,105,110,103,32,111,102,32,116,104,101,32,119,111,114,108,100,
44,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,62,32,66,117,116,32,119,101,32,105,110,32,105,116,32,115,104,97,
108,108,32,98,101,32,114,101,109,101,109,98,101,114,101,100,45,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,62,32,87,101,32,102,101,119,44,32,119,101,32,104,97,112,112,121,32,
102,101,119,44,32,119,101,32,98,97,110,100,32,111,102,32,98,114,111,116,104,101,
114,115,59,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,62,32,70,111,114,32,104,101,32,116,111,45,100,97,121,32,116,
104,97,116,32,115,104,101,100,115,32,104,105,115,32,98,108,111,111,100,32,119,105,
116,104,32,109,101,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,83,104,97,108,108,32,98,101,32,109,121,32,98,
114,111,116,104,101,114,59,32,98,101,32,104,101,32,110,101,39,101,114,32,115,111,
32,118,105,108,101,44,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,84,104,105,115,32,100,97,121,32,115,104,
97,108,108,32,103,101,110,116,108,101,32,104,105,115,32,99,111,110,100,105,116,
105,111,110,59,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,65,110,100,32,103,101,110,116,108,101,
109,101,110,32,105,110,32,69,110,103,108,97,110,100,32,110,111,119,45,97,45,98,
101,100,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,83,104,97,108,108,32,116,104,105,110,107,
32,116,104,101,109,115,101,108,118,101,115,32,97,99,99,117,114,115,39,100,32,116,
104,101,121,32,119,101,114,101,32,110,111,116,32,104,101,114,101,44,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,60,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,62,32,65,110,100,32,
104,111,108,100,32,116,104,101,105,114,32,109,97,110,104,111,111,100,115,32,99,
104,101,97,112,32,119,104,105,108,101,115,32,97,110,121,32,115,112,101,97,107,115,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,60,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
62,32,84,104,97,116,32,102,111,117,103,104,116,32,119,105,116,104,32,117,115,32,
117,112,111,110,32,83,97,105,110,116,32,67,114,105,115,112,105,110,39,115,32,100,
97,121,46,32,32,32,32,32,32,32,32,83,104,97,107,101,115,112,101,97,114,101,44,32,
72,101,110,114,121,32,86,44,32,65,99,116,32,73,86,44,32,83,99,101,110,101,32,51,
60,0,others=>0);

signal addr1: integer range 0 to 8191; -- address for memory port 1 (display side)
signal addr2: integer range 0 to 8191; -- address for memory port 2 (serial side)
type state_type is (idle, scrolling, clearing);
signal nxt,cur: state_type;
signal we, seq_comp, seq_go: std_logic;
signal seq_col: integer range 0 to 92;
signal seq_row: integer range 0 to 47;
signal row: std_logic_vector(5 downto 0);
signal col: std_logic_vector(6 downto 0);
signal data_in, data_out: std_logic_vector(6 downto 0);

  
begin

process(clk)
begin
	if rising_edge(clk) then
		cur <= nxt;
	end if;
end process;

--Controller
process(cur, seq_comp, scroll, clear)
begin
we <= '0';
seq_go <= '0';
	case cur is
		when idle => 
			seq_go <= scroll or clear;
			we <= writec;
			if clear = '1' then
				nxt <= clearing;
			elsif scroll = '1' then
				nxt <= scrolling;
			else
				nxt <= idle;
			end if;
		when clearing =>
			we <= '1';
			if seq_comp = '0' then
				nxt <= clearing;
			else
				nxt <= idle;
			end if;
		when scrolling =>
			we <= '1';
			if seq_comp = '0' then
				nxt <= scrolling;
			else
				nxt <= idle;
			end if;
	end case;
end process;

--seq_row 0 -> 47, seq_col 0 -> 92
process(clk) 
begin
	if rising_edge(clk) then
		if seq_go = '1' then
			seq_col <= 92;
			seq_row <= 47;
		elsif seq_row /= 0 then
			seq_row <= seq_row - 1;
		elsif seq_col /= 0 then
			seq_row <= 47;
			seq_col <= seq_col - 1;
		end if;
	end if;
end process;

--Sequence Complete
seq_comp <= '1' when seq_row = 0 and seq_col = 0 else '0';
-- Row and Col Mux's
row <= row2 when cur = idle else std_logic_vector(to_unsigned(seq_row,row'length));
col <= col2 when cur = idle else std_logic_vector(to_unsigned(seq_col,col'length));
-- Ascii2 Mux
data_in <= "0000000" when cur = clearing or (cur = scrolling and seq_row = 47) else data_out when cur = scrolling else in2;

--   model output (display side) of character memory - use block memory
  addr1 <= to_integer(unsigned(row1&col1));
  process (clk)
  begin
    if rising_edge(clk) then
      out1 <= std_logic_vector(to_unsigned(char_ram(addr1),7));
    end if;
  end process;
  
  -- model input (serial side) of character memory - use block memory
  addr2 <= to_integer(unsigned(row & col));
  process (clk)
  begin
    if rising_edge(clk) then
      if we = '1' then
        char_ram(addr2)<=to_integer(unsigned(data_in));
      end if;
      data_out <= std_logic_vector(to_unsigned(char_ram(addr2),7));
    end if;
  end process;

end behavioral;
