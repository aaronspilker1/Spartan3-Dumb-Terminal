----------------------------------------------------------------------------------
-- Company: Weber State
-- Engineer: Aaron Spilker
-- Module Name:    char_gen - Behavioral 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity chargen is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           hstart : in  STD_LOGIC;
           vga_row : in  STD_LOGIC_VECTOR (9 downto 0);
			  ascii: in STD_LOGIC_VECTOR (6 downto 0);
			  row_addr: out STD_LOGIC_VECTOR (5 downto 0);
			  col_addr: out STD_LOGIC_VECTOR (6 downto 0);
           pix : out  STD_LOGIC);
end chargen;

architecture Behavioral of chargen is
  -- 11x16 font
  -- each character has 16 words, each of which are 11 bits. The array below is actually 12 bits wide to
  -- facilitate initialization with the X"hhh" notation. Ignore the most significant bit. There are 128
  -- characters in all, but the first 32 are unprintable control characters. All those characters render
  -- as blanks. The same is true for character 127 (7F). The first word of any character represents the
  -- top row of pixels in that character. The sixteenth word represents the bottom row of pixels.
 type font_rom_type is array (0 to 2047) of unsigned(11 downto 0);
 
 constant font_rom: font_rom_type := (
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- NUL
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- SOH
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- STX
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- ETX
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- EOT
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- ENQ
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- ACK
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- BEL
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- BS
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- TAB
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- LF
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- VT
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- FF
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- CR
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- SO
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- SI
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- DLE
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- DC1
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- DC2
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- DC3
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- DC4
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- NAK
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- SYN
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- ETB
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- CAN
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- EM
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- SUB
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- ESC
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- FS
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- GS
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- RS
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- US
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- space
    X"000",X"000",X"000",X"040",X"040",X"040",X"040",X"040",X"040",X"000",X"000",X"040",X"000",X"000",X"000",X"000", -- !
    X"000",X"000",X"000",X"090",X"090",X"090",X"090",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- "
    X"000",X"000",X"090",X"090",X"090",X"3fc",X"090",X"090",X"3fc",X"090",X"090",X"090",X"000",X"000",X"000",X"000", -- #
    X"000",X"040",X"040",X"0f0",X"110",X"100",X"180",X"060",X"018",X"008",X"108",X"1f0",X"040",X"040",X"000",X"000", -- $
    X"000",X"000",X"000",X"1c0",X"220",X"224",X"1d8",X"060",X"1b8",X"244",X"044",X"038",X"000",X"000",X"000",X"000", -- %
    X"000",X"000",X"000",X"0c0",X"120",X"100",X"080",X"1d8",X"250",X"230",X"230",X"1dc",X"000",X"000",X"000",X"000", -- &
    X"000",X"000",X"000",X"040",X"040",X"040",X"040",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- '
    X"000",X"000",X"000",X"010",X"020",X"020",X"040",X"040",X"040",X"040",X"040",X"040",X"020",X"020",X"010",X"000", -- (
    X"000",X"000",X"000",X"100",X"080",X"080",X"040",X"040",X"040",X"040",X"040",X"040",X"080",X"080",X"100",X"000", -- )
    X"000",X"000",X"088",X"050",X"020",X"1fc",X"020",X"050",X"088",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- *
    X"000",X"000",X"000",X"000",X"020",X"020",X"020",X"1fc",X"020",X"020",X"020",X"000",X"000",X"000",X"000",X"000", -- +
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"060",X"040",X"040",X"080",X"000",X"000", -- ,
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"1f8",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- -
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"070",X"070",X"000",X"000",X"000",X"000", -- .
    X"000",X"000",X"008",X"010",X"010",X"020",X"020",X"040",X"040",X"040",X"080",X"080",X"100",X"000",X"000",X"000", -- /
    X"000",X"000",X"0f0",X"108",X"108",X"108",X"108",X"108",X"108",X"108",X"108",X"0f0",X"000",X"000",X"000",X"000", -- 0
    X"000",X"000",X"0c0",X"140",X"240",X"040",X"040",X"040",X"040",X"040",X"040",X"3f8",X"000",X"000",X"000",X"000", -- 1
    X"000",X"000",X"1e0",X"210",X"010",X"010",X"010",X"020",X"040",X"080",X"110",X"3f0",X"000",X"000",X"000",X"000", -- 2
    X"000",X"000",X"1e0",X"210",X"010",X"010",X"0e0",X"010",X"010",X"010",X"210",X"1e0",X"000",X"000",X"000",X"000", -- 3
    X"000",X"000",X"030",X"050",X"050",X"090",X"110",X"110",X"210",X"3f8",X"010",X"078",X"000",X"000",X"000",X"000", -- 4
    X"000",X"000",X"1f0",X"100",X"100",X"100",X"1f0",X"108",X"008",X"008",X"208",X"1f0",X"000",X"000",X"000",X"000", -- 5
    X"000",X"000",X"078",X"080",X"080",X"100",X"170",X"188",X"108",X"108",X"088",X"070",X"000",X"000",X"000",X"000", -- 6
    X"000",X"000",X"3f0",X"210",X"020",X"020",X"020",X"040",X"040",X"040",X"080",X"080",X"000",X"000",X"000",X"000", -- 7
    X"000",X"000",X"0f0",X"108",X"108",X"108",X"0f0",X"090",X"108",X"108",X"108",X"0f0",X"000",X"000",X"000",X"000", -- 8
    X"000",X"000",X"0e0",X"110",X"108",X"108",X"118",X"0e8",X"008",X"010",X"010",X"1e0",X"000",X"000",X"000",X"000", -- 9
    X"000",X"000",X"000",X"000",X"000",X"070",X"070",X"000",X"000",X"000",X"070",X"070",X"000",X"000",X"000",X"000", -- :
    X"000",X"000",X"000",X"000",X"000",X"070",X"070",X"000",X"000",X"000",X"070",X"060",X"0c0",X"0c0",X"000",X"000", -- ;
    X"000",X"000",X"000",X"000",X"00c",X"030",X"0c0",X"300",X"0c0",X"030",X"00c",X"000",X"000",X"000",X"000",X"000", -- <
    X"000",X"000",X"000",X"000",X"000",X"000",X"1fc",X"000",X"000",X"1fc",X"000",X"000",X"000",X"000",X"000",X"000", -- =
    X"000",X"000",X"000",X"000",X"300",X"0c0",X"030",X"00c",X"030",X"0c0",X"300",X"000",X"000",X"000",X"000",X"000", -- >
    X"000",X"000",X"000",X"0f0",X"108",X"008",X"010",X"020",X"020",X"000",X"020",X"020",X"000",X"000",X"000",X"000", -- ?
    X"000",X"000",X"0e0",X"110",X"210",X"270",X"2d0",X"290",X"290",X"2f8",X"110",X"0e0",X"000",X"000",X"000",X"000", -- @
    X"000",X"000",X"000",X"0f0",X"030",X"030",X"048",X"048",X"0fc",X"084",X"084",X"3ce",X"000",X"000",X"000",X"000", -- A
    X"000",X"000",X"000",X"3f0",X"108",X"108",X"108",X"1f0",X"108",X"104",X"104",X"3f8",X"000",X"000",X"000",X"000", -- B
    X"000",X"000",X"000",X"0f4",X"10c",X"204",X"200",X"200",X"200",X"200",X"104",X"0f8",X"000",X"000",X"000",X"000", -- C
    X"000",X"000",X"000",X"3f0",X"108",X"104",X"104",X"104",X"104",X"104",X"108",X"3f0",X"000",X"000",X"000",X"000", -- D
    X"000",X"000",X"000",X"3fc",X"104",X"104",X"110",X"1f0",X"110",X"104",X"104",X"3fc",X"000",X"000",X"000",X"000", -- E
    X"000",X"000",X"000",X"3f8",X"108",X"108",X"120",X"1e0",X"120",X"100",X"100",X"380",X"000",X"000",X"000",X"000", -- F
    X"000",X"000",X"000",X"0f4",X"10c",X"204",X"200",X"200",X"21e",X"204",X"104",X"0fc",X"000",X"000",X"000",X"000", -- G
    X"000",X"000",X"000",X"39c",X"108",X"108",X"108",X"1f8",X"108",X"108",X"108",X"39c",X"000",X"000",X"000",X"000", -- H
    X"000",X"000",X"000",X"1f0",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"1f0",X"000",X"000",X"000",X"000", -- I
    X"000",X"000",X"000",X"0f8",X"010",X"010",X"010",X"210",X"210",X"210",X"310",X"1e0",X"000",X"000",X"000",X"000", -- J
    X"000",X"000",X"000",X"3bc",X"110",X"120",X"140",X"1c0",X"120",X"110",X"108",X"39e",X"000",X"000",X"000",X"000", -- K
    X"000",X"000",X"000",X"380",X"100",X"100",X"100",X"100",X"108",X"108",X"108",X"3f8",X"000",X"000",X"000",X"000", -- L
    X"000",X"000",X"000",X"71c",X"318",X"2a8",X"2a8",X"2a8",X"248",X"248",X"208",X"79c",X"000",X"000",X"000",X"000", -- M
    X"000",X"000",X"000",X"73c",X"308",X"288",X"288",X"248",X"228",X"228",X"218",X"798",X"000",X"000",X"000",X"000", -- N
    X"000",X"000",X"000",X"0f0",X"108",X"204",X"204",X"204",X"204",X"204",X"108",X"0f0",X"000",X"000",X"000",X"000", -- O
    X"000",X"000",X"000",X"1f8",X"084",X"084",X"084",X"084",X"0f8",X"080",X"080",X"1e0",X"000",X"000",X"000",X"000", -- P
    X"000",X"000",X"000",X"0f0",X"108",X"204",X"204",X"204",X"204",X"30c",X"108",X"0f0",X"060",X"09c",X"000",X"000", -- Q
    X"000",X"000",X"000",X"3f0",X"108",X"108",X"108",X"1f0",X"120",X"110",X"108",X"38c",X"000",X"000",X"000",X"000", -- R
    X"000",X"000",X"000",X"0f4",X"10c",X"104",X"100",X"0f8",X"004",X"104",X"184",X"178",X"000",X"000",X"000",X"000", -- S
    X"000",X"000",X"000",X"3f8",X"248",X"248",X"040",X"040",X"040",X"040",X"040",X"0e0",X"000",X"000",X"000",X"000", -- T
    X"000",X"000",X"000",X"73c",X"208",X"208",X"208",X"208",X"208",X"208",X"110",X"0e0",X"000",X"000",X"000",X"000", -- U
    X"000",X"000",X"000",X"39c",X"108",X"108",X"108",X"090",X"090",X"090",X"060",X"060",X"000",X"000",X"000",X"000", -- V
    X"000",X"000",X"000",X"38e",X"104",X"124",X"154",X"154",X"154",X"0d8",X"088",X"088",X"000",X"000",X"000",X"000", -- W
    X"000",X"000",X"000",X"38e",X"104",X"088",X"050",X"020",X"050",X"088",X"104",X"38e",X"000",X"000",X"000",X"000", -- X
    X"000",X"000",X"000",X"71c",X"208",X"110",X"0a0",X"0a0",X"040",X"040",X"040",X"0e0",X"000",X"000",X"000",X"000", -- Y
    X"000",X"000",X"000",X"3f8",X"208",X"210",X"020",X"040",X"080",X"108",X"208",X"3f8",X"000",X"000",X"000",X"000", -- Z
    X"000",X"000",X"000",X"070",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"070",X"000", -- [
    X"000",X"000",X"000",X"100",X"080",X"080",X"040",X"040",X"020",X"020",X"010",X"010",X"008",X"000",X"000",X"000", -- \
    X"000",X"000",X"000",X"1c0",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"1c0",X"000", -- ]
    X"000",X"000",X"000",X"020",X"050",X"088",X"104",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- ^
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"7ff",X"000", -- _
    X"000",X"180",X"0c0",X"040",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- `
    X"000",X"000",X"000",X"000",X"000",X"0f0",X"108",X"008",X"1f8",X"208",X"218",X"1ec",X"000",X"000",X"000",X"000", -- a
    X"000",X"000",X"380",X"080",X"080",X"0b8",X"0c4",X"082",X"082",X"082",X"0c4",X"1b8",X"000",X"000",X"000",X"000", -- b
    X"000",X"000",X"000",X"000",X"000",X"074",X"08c",X"104",X"100",X"100",X"084",X"078",X"000",X"000",X"000",X"000", -- c
    X"000",X"000",X"038",X"008",X"008",X"0e8",X"118",X"208",X"208",X"208",X"118",X"0ec",X"000",X"000",X"000",X"000", -- d
    X"000",X"000",X"000",X"000",X"000",X"1f8",X"204",X"204",X"3fc",X"200",X"204",X"1f8",X"000",X"000",X"000",X"000", -- e
    X"000",X"000",X"03c",X"040",X"040",X"1fc",X"040",X"040",X"040",X"040",X"040",X"0fc",X"000",X"000",X"000",X"000", -- f
    X"000",X"000",X"000",X"000",X"000",X"0ec",X"118",X"208",X"208",X"208",X"118",X"0e8",X"008",X"008",X"1f0",X"000", -- g
    X"000",X"000",X"380",X"080",X"080",X"0b8",X"0c4",X"084",X"084",X"084",X"084",X"1ce",X"000",X"000",X"000",X"000", -- h
    X"000",X"020",X"020",X"000",X"000",X"060",X"020",X"020",X"020",X"020",X"020",X"1fc",X"000",X"000",X"000",X"000", -- i
    X"000",X"008",X"008",X"000",X"000",X"0f8",X"008",X"008",X"008",X"008",X"008",X"008",X"008",X"018",X"0f0",X"000", -- j
    X"000",X"000",X"380",X"080",X"080",X"09c",X"090",X"0a0",X"0c0",X"0b0",X"088",X"19e",X"000",X"000",X"000",X"000", -- k
    X"000",X"000",X"1e0",X"020",X"020",X"020",X"020",X"020",X"020",X"020",X"020",X"1fc",X"000",X"000",X"000",X"000", -- l
    X"000",X"000",X"000",X"000",X"000",X"3d8",X"124",X"124",X"124",X"124",X"124",X"3b6",X"000",X"000",X"000",X"000", -- m
    X"000",X"000",X"000",X"000",X"000",X"1b8",X"0c4",X"084",X"084",X"084",X"084",X"1ce",X"000",X"000",X"000",X"000", -- n
    X"000",X"000",X"000",X"000",X"000",X"0f0",X"108",X"204",X"204",X"204",X"108",X"0f0",X"000",X"000",X"000",X"000", -- o
    X"000",X"000",X"000",X"000",X"000",X"370",X"188",X"104",X"104",X"104",X"188",X"170",X"100",X"100",X"3c0",X"000", -- p
    X"000",X"000",X"000",X"000",X"000",X"0ec",X"118",X"208",X"208",X"208",X"118",X"0e8",X"008",X"008",X"03c",X"000", -- q
    X"000",X"000",X"000",X"000",X"000",X"19c",X"0e0",X"080",X"080",X"080",X"080",X"1f0",X"000",X"000",X"000",X"000", -- r
    X"000",X"000",X"000",X"000",X"000",X"0fc",X"104",X"100",X"0f8",X"004",X"104",X"1f8",X"000",X"000",X"000",X"000", -- s
    X"000",X"000",X"000",X"080",X"080",X"1f8",X"080",X"080",X"080",X"080",X"084",X"078",X"000",X"000",X"000",X"000", -- t
    X"000",X"000",X"000",X"000",X"000",X"318",X"108",X"108",X"108",X"108",X"118",X"0ec",X"000",X"000",X"000",X"000", -- u
    X"000",X"000",X"000",X"000",X"000",X"3ce",X"084",X"084",X"048",X"048",X"030",X"030",X"000",X"000",X"000",X"000", -- v
    X"000",X"000",X"000",X"000",X"000",X"38e",X"202",X"124",X"154",X"154",X"0d8",X"0d8",X"000",X"000",X"000",X"000", -- w
    X"000",X"000",X"000",X"000",X"000",X"39c",X"108",X"090",X"060",X"090",X"108",X"39c",X"000",X"000",X"000",X"000", -- x
    X"000",X"000",X"000",X"000",X"000",X"70e",X"108",X"108",X"090",X"090",X"060",X"020",X"040",X"080",X"3e0",X"000", -- y
    X"000",X"000",X"000",X"000",X"000",X"1f8",X"110",X"020",X"040",X"040",X"088",X"1f8",X"000",X"000",X"000",X"000", -- z
    X"000",X"000",X"000",X"030",X"040",X"040",X"040",X"040",X"040",X"080",X"040",X"040",X"040",X"040",X"030",X"000", -- {
    X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040",X"040", -- |
    X"000",X"000",X"000",X"0c0",X"020",X"020",X"020",X"020",X"020",X"010",X"020",X"020",X"020",X"020",X"0c0",X"000", -- }
    X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"1c4",X"238",X"000",X"000",X"000",X"000",X"000",X"000",X"000", -- ~
    X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF",X"FFF"); -- DEL

signal count: integer range 0 to 10;
signal col: integer range 0 to 93;
signal load: std_logic;
signal font: std_logic_vector(11 downto 0);
signal to_font: std_logic_vector(10 downto 0);

begin
col_addr <= std_logic_vector(to_unsigned(col,col_addr'length));
row_addr <= vga_row(9 downto 4); 
to_font <= ascii & vga_row(3 downto 0);
load <= '1' when hstart = '1' or count = 10 else '0';

--Column Counter (0-10)
process(clk)
begin
	if rising_edge(clk) then
		if hstart = '1' or count = 10 then
			count <= 0;
		else
			count <= count + 1;
		end if;
	end if;
end process;

--Column Counter (0-92)
process(clk,reset)
begin 
	if reset = '1' then
		col <= 0;
	elsif rising_edge(clk) then
		if load = '1' then
			if col = 93 then
				col <= 0;
			elsif col /= 0 then
				col <= col + 1;
			elsif hstart = '1' then
				col <= 1;
			end if;
		end if;
	end if;
end process;

--every 11 clock cycles shift Q10 to pixel out.
pix <= font(10);

process(clk)
begin
	if rising_edge(clk) then
		if load = '1' then
			font <= std_logic_vector(font_rom(to_integer(unsigned(to_font)))); -- font for shift register 
		else
			font <= font(10 downto 0) & '0';
		end if;
	end if;
end process;

end Behavioral;
